0
2 2 2 2 2 r 0 2 h 0 T 2 T
1 2 2 2 2 r h 4 T
2 2 2 2 2 r h 6 T
4 3 3 3 3 r h 8 T
2 3 1 12 4 2 4 12 3 9 3 6 2 4 1 10 2 2 0 5 4 5 0 8 0 8 1 8 3 4 1 12 2 2 5 7 0 11
