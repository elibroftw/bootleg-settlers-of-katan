0
2 2 2 2 2 r 7 15 h 0 T 2 T 4 T
0 0 0 0 0 r h
0 0 0 0 0 r h
0 0 0 0 0 r h
2 3 1 12 4 2 4 12 3 9 3 6 2 4 1 10 2 2 0 5 4 5 0 8 0 8 1 8 3 4 1 12 2 2 5 7 0 11
