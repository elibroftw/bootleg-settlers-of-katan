0
2 2 2 2 2 r 0 2 h 0 T 2 T
1 2 2 2 2 r h 4 T
2 2 2 2 2 r h 6 T
4 3 3 3 3 r h 8 T
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
